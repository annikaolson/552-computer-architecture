module decode_stage();

// decoding the instructions

endmodule