module write_back_stage();

// reg file write (assert signals)

endmodule