module memory_stage();

// read to or write from memory
// pc = target if beq

endmodule