module fetch_stage();


// instr = mem[pc]
// new pc set up

endmodule