module execute_stage();

// aluout = rs op rt 
// branch target gets computed


endmodule